// ----------------------------------------------------------------------------
// arty_test_pkg.sv
//
// 9/1/2025 D. Hawkins (dwh@caltech.edu)
//
// Digilent Arty test package.
//
// ----------------------------------------------------------------------------

`timescale 1ps / 1ps

package arty_test_pkg;

	// ------------------------------------------------------------------------
	// Packages
	// ------------------------------------------------------------------------
	//
	// Vivado AXI4-MM Verification IP
	import axi_vip_pkg::*;

	// Custom packages
	import aximm_memory_pkg::*;

	// ----------------------------------------------------------------------------
	// Test Class
	// ----------------------------------------------------------------------------
	//
	`include "arty_test.svh"

endpackage
