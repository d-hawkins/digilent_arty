// ----------------------------------------------------------------------------
// aximm_gpio_pkg.sv
//
// 9/1/2025 D. W. Hawkins (dwh@caltech.edu)
//
// AXI-MM GPIO test package.
//
// ----------------------------------------------------------------------------

package aximm_gpio_pkg;

	// ------------------------------------------------------------------------
	// Packages
	// ------------------------------------------------------------------------
	//
	import aximm_base_pkg::*;

	// ------------------------------------------------------------------------
	// AXI4-MM GPIO Control/Status
	// ------------------------------------------------------------------------
	//
	class aximm_gpio #(type AXIMM) extends aximm_base #(AXIMM);

		// --------------------------------------------------------------------
		// Member Variables
		// --------------------------------------------------------------------
		//
		// GPIO base address
		int m_addr;

		// --------------------------------------------------------------------
		// Member Functions
		// --------------------------------------------------------------------
		//
		// Constructor
		function new(
			AXIMM axi,
			int   base_addr
		);
			// Baseclass constructor
			super.new(axi);

			// Extended class
			m_addr = base_addr;
		endfunction

		// --------------------------------------------------------------------
		// Member Tasks
		// --------------------------------------------------------------------
		//
		// --------------------------------------------------------------------
		// Control Write
		// --------------------------------------------------------------------
		//
		task control_write (
			input int unsigned data
		);
			axi_write_single(m_addr+0, data);
		endtask

		// --------------------------------------------------------------------
		// Control Read
		// --------------------------------------------------------------------
		//
		task control_read (
			output int unsigned data
		);
			axi_read_single(m_addr+0, data);
		endtask

		// --------------------------------------------------------------------
		// Status Read
		// --------------------------------------------------------------------
		//
		task status_read (
			output int unsigned data
		);
			axi_read_single(m_addr+8, data);
		endtask
	endclass
endpackage

